//-------------------------------------------------------------------------------
//  FEUP / MEEC - Digital Systems Design 2023/2024
//
//  jca@fe.up.pt, Nov 2023
// 
// 	This Verilog code is property of University of Porto
// 	Its utilization beyond the scope of the course Digital Systems Design
// 	(Projeto de Sistemas Digitais) of the Master in Electrical 
// 	and Computer Engineering requires explicit authorization from the author.
// 
//-------------------------------------------------------------------------------
`timescale 1ns/100ps
module cpxdiv_tb;

// Signals to connect to your cpxdiv module:
reg clock;
reg reset;
reg run;
reg [15:0] ReA;
reg [15:0] ImA;
reg [15:0] ReB;
reg [15:0] ImB;
wire [31:0] ReY;
wire [31:0] ImY;
wire busy;


// Instantiate the circuit under verification
// Note this is "golden" simulation model, you must change it to your module:
cpxdiv3  mycpxdiv(
         .clock( clock ),
         .reset( reset ),
         .run( run ),
         .ReA( ReA ),
         .ImA( ImA ),
         .ReB( ReB ),
         .ImB( ImB ),
         .ReY( ReY ),
         .ImY( ImY ),
         .busy( busy )
             );



// The good expected results generated by "golden" tasks:
reg [31:0] GoldenReY;
reg [31:0] GoldenImY;

// The errors: obtained - expected
reg [31:0] err_Re = 0, err_Im = 0;

// Float operands:
real fReA, fImA, fReB, fImB, fReY, fImY;

// Set FULL_DEBUG to 1 to print intermediate results of the fixed-point calculation
// Set PRINT_RESULTS to 1 to print all results
integer FULL_DEBUG      = 0,
        PRINT_RESULTS   = 1;


// Set initial values, generate the clock signal:
initial
begin
  clock = 0;
  reset = 0;
  ReA = 0;
  ImA = 0;
  ReB = 0;
  ImB = 0;
  run = 0;
  #2
  // free running clock signal:
  forever #2.5 clock = ~clock;
end

// Simple reset, one clock period aligned with the negedge of the clock:
initial
begin
  #1
  #200
  @(negedge clock);
  reset = 1;
  @(negedge clock);
  reset = 0;
end


// Main verification program
initial
begin

  FULL_DEBUG = 0;
  PRINT_RESULTS = 1;
  
  // How to use the verification tasks:

  // First examples calculate and print various complex divisions
  // This is just to test the verification tasks:
  
  // Set float operands in the range [-128.0, +127.0]:
  fReA = 123.45;    fImA = 65.27;
  fReB = 56.71;     fImB = 12.345;
  
  // Calculate the complex division and print results obtained by 3 different processes:
  // i)   using the float input variables and float arithmetic operation (full Verilog precision)
  // ii)  using the fixed-point input variables (converted to float) and float arithmetic
  // iii) using the fixed-point input variables (as integers) and fixed-point arithmetic
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );


  // Experiment with some other cases, with negative and positive operands:
  fReA = -124.45;   fImA = 65.27;
  fReB = 56.71;     fImB = 12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = -102.76;    fImA = 65.27;
  fReB = 36.79;      fImB = -12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = 123.45;    fImA = -65.27;
  fReB = 56.71;     fImB = -12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = 123.45;    fImA = -65.27;
  fReB = -0.71;     fImB = -1.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = 18.45;    fImA = -65.27;
  fReB = 5.25;     fImB = -12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = 18.45;    fImA = -65.27;
  fReB = -5.25;     fImB = -12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = -18.45;    fImA = -65.27;
  fReB = -5.25;     fImB = -12.345;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );

  fReA = 123.45;    fImA = -65.27;
  fReB = 2.01;     fImB = -0.25;
  golden_cpxdiv( fReA, fImA, fReB, fImB, fReY, fImY );


 
  //----------------------------------------------------------------------------
  // How to build your testbench:
  
  // Your circuit is connected to the registers ReA, ImA, ReB and ImB
  // and the outputs are connected to ReY[31:0] and ImY[31:0]
  // one verification can be implementes as:
  
  #1
  @(negedge reset) // Block until reset is released
  repeat (10)
    @(negedge clock); // Wait some clock cycles before starting the operation
	
  // Set float operands:
  fReA = 123.45;    fImA = -65.27;  fReB = 2.01;     fImB = -0.25;
  
  // Convert float operands f* to 16-bit fixed-point, with 8-fractional bit:
  // The registers ReA, ImA, ReB and ImB (16-bit signed integers) are the inputs
  // to apply to your complex divisor:
  ReA = fReA * 256;  ImA = fImA * 256;  ReB = fReB * 256;  ImB = fImB * 256;
  
  // Your complex divisor outputs two 32-bit signed integers ReY and ImY, representing 
  // the real and imaginary parts of the result. To obtain the expected values for ReY and ImY
  // (the "golden" values) call the task golden_cpxdiv_fxpoint( ReA, ImA, ReB, ImB, GoldenReY, GoldenImY ); 
  // NOTE this is also done within the task golden_cpxdiv( ) used above:
  golden_cpxdiv_fxpoint( ReA, ImA, ReB, ImB, GoldenReY, GoldenImY );
  
  // Start your module and wait for the end of the calculation process:
  
 
  @(negedge clock); // Synchronize with the negative edge of the clock signal
  run = 1;   // Start the complex divider, set run to 1 for one clock period
  @(negedge clock); 
  run = 0;
  @(negedge clock); 
  while ( busy == 1 ) @(negedge clock);  // Wait for busy low. When busy is low the results should be at the output ports
  
  // Errors:
  err_Re = ReY - GoldenReY;
  err_Im = ImY - GoldenImY;
  
  // Compare the results generated by your circuit in the wires ReY and ImY
  // with the expected golden results computed by task golden_cpxdiv_fxpoint( ) in GoldenReY and GoldenImY:
  if ( ReY !== GoldenReY || ImY !== GoldenImY )
  begin
    // do something when an error is found !
	// Print as 32-bit signed integers:
	if (PRINT_RESULTS) $write("ERROR: Expected (as integers): %d + j %d, obtained %d + j %d\n", 
	                                   $signed(GoldenReY), $signed(GoldenImY), $signed(ReY), $signed(ImY) );
									   
	// And/or print as 32-bit fixed-point with 16 fractional bits:
	if (PRINT_RESULTS) $write("ERROR: Expected (as floats)  : %1.8f + j %1.8f, obtained %1.8f + j %1.8f\n", 
	                                   $signed(GoldenReY)/65536.0, $signed(GoldenImY)/65536.0,
									   $signed(ReY)/65536.0, $signed(ImY)/65536.0 );
	
	$stop; // Stop if an error is found
  end
  

  
  $stop;
  
end



//--------------------------------------------------------------------
// Check range of operands, calculate and print the complex division for:
// i)  using the float input variables and float arithmetic operation (full Verilog precision)
// ii) using the fixed-point input variables (converted to float) and float arithmetic
// iii)using the fixed-point input variables (as integers) and fixed-point arithmetic
task golden_cpxdiv( 
                    input  real fReA,
					input  real fImA,
					input  real fReB,
					input  real fImB,
					output real fReY,
					output real fImY
					);
					
reg [15:0] ReA;
reg [15:0] ImA;
reg [15:0] ReB;
reg [15:0] ImB;
reg [31:0] ReY;
reg [31:0] ImY;

// Float operands, fractional part truncated to 8 bits:
real fpReA, fpImA, fpReB, fpImB;
// Float results:
real fpReY, fpImY;					
begin					
	
  if (PRINT_RESULTS) $write("----------------------------------------------------------------------------------------------\n");
	
  // Test the range of the operands:
  if ( fReA > 127.0 || fReA < -128.0 ||
       fReB > 127.0 || fReB < -128.0 ||
	   fImA > 127.0 || fImA < -128.0 ||
	   fImB > 127.0 || fImB < -128.0 
	   )
  begin
    // Out of range, print error and return
	if (PRINT_RESULTS) $write("######################################################################\n");
    if (PRINT_RESULTS) $write( "Operands out of range: A = (%1.8f + j %1.8f )\n", fReA, fImA );
    if (PRINT_RESULTS) $write( "                       B = (%1.8f + j %1.8f )\n", fReB, fImB );
	if (PRINT_RESULTS) $write( "The real and imaginary parts must be in [-128.0, +127.0]\n");
	if (PRINT_RESULTS) $write("######################################################################\n");
  end
  else
  begin
  
	// Calculate the complex division with float input data using full precision float arithmetic:					
    golden_cpxdiv_float( fReA, fImA, fReB, fImB, fReY, fImY );
    if (PRINT_RESULTS) $write("Float full precision        : (%1.8f + j %1.8f ) / (%1.8f + j %1.8f ) = %1.8f + j %1.8f \n",
                                            fReA, fImA, fReB, fImB, fReY, fImY );   
    
    // Convert float input operands to 16-bit integers:
    ReA = fReA * 256;
    ImA = fImA * 256;
    ReB = fReB * 256;
    ImB = fImB * 256;
	
	// Convert back to float, fractional is part truncated to 8 bits
    fpReA = $signed(ReA) / 256.0;
    fpImA = $signed(ImA) / 256.0;
    fpReB = $signed(ReB) / 256.0;
    fpImB = $signed(ImB) / 256.0;
	
	// Calculate the complex division with the fixed-point input data, truncated to 8 fractional bits
	// using full precision float arithmetic:
    golden_cpxdiv_float( fpReA, fpImA, fpReB, fpImB, fpReY, fpImY );
    if (PRINT_RESULTS) $write("Fixed-point data, float calc: (%1.8f + j %1.8f ) / (%1.8f + j %1.8f ) = %1.8f + j %1.8f \n",
                                            fpReA, fpImA, fpReB, fpImB, fpReY, fpImY );   
    
	// Calculate the complex division with the fixed-point input data, truncated to 8 fractional bits
	// using fixed-point precision arithmetic, as specified for the project:
    golden_cpxdiv_fxpoint( ReA, ImA, ReB, ImB, ReY, ImY );	  
    if (PRINT_RESULTS) $write("Fixed-point data and calc   : (%1.8f + j %1.8f ) / (%1.8f + j %1.8f ) = %1.8f + j %1.8f \n",
                                            fpReA, fpImA, fpReB, fpImB, $signed(ReY)/65536.0, $signed(ImY)/65536.0 );
  end
	  
end
endtask		



//--------------------------------------------------------------------
// Complex division with float data calculated in full float precision
task golden_cpxdiv_float(
                        input real ReA,
					    input real ImA,
					    input real ReB,
					    input real ImB,
						output real ReY,
						output real ImY
					   );
begin
  ReY = ( ReA * ReB + ImA * ImB ) / ( ReB * ReB + ImB * ImB );
  ImY = ( ReB * ImA - ReA * ImB ) / ( ReB * ReB + ImB * ImB );
end
endtask


//--------------------------------------------------------------------
// Complex division with fixed-point data and calculated in fixed-point:
task golden_cpxdiv_fxpoint(
                        input [15:0] ReA,
					    input [15:0] ImA,
					    input [15:0] ReB,
					    input [15:0] ImB,
						output [31:0] ReY,
						output [31:0] ImY
					   );
reg signed [31:0] P1, P2, P3, P4, P5, P6;
reg signed [31:0] NumeR, NumeI;
reg        [31:0] Denom;				   
begin
  P1 = fxpmult( ReA, ReB );
  P2 = fxpmult( ImA, ImB );
  P3 = fxpmult( ReB, ImA );
  P4 = fxpmult( ReA, ImB );
  P5 = fxpmult( ReB, ReB );
  P6 = fxpmult( ImB, ImB );
  
  NumeR = P1 + P2; // ( ReA * ReB + ImA * ImB )
  NumeI = P3 - P4; // ( ReB * ImA - ReA * ImB )
  Denom = P5 + P6; // ( ReB * ReB + ImB * ImB )

  ReY = fxpdiv( NumeR, Denom[31:16] );
  ImY = fxpdiv( NumeI, Denom[31:16] );
  
  if ( FULL_DEBUG )
  begin
    if (PRINT_RESULTS) $write("ReA * ReB = %d (%1.8f)\n", P1, P1/65536.0 );
    if (PRINT_RESULTS) $write("ImA * ImB = %d (%1.8f)\n", P2, P2/65536.0 );
    if (PRINT_RESULTS) $write("ReB * ImA = %d (%1.8f)\n", P3, P3/65536.0 );
    if (PRINT_RESULTS) $write("ReA * ImB = %d (%1.8f)\n", P4, P4/65536.0 );
    if (PRINT_RESULTS) $write("ReB * ImB = %d (%1.8f)\n", P5, P5/65536.0 );
    if (PRINT_RESULTS) $write("ImB * ImB = %d (%1.8f)\n", P6, P6/65536.0 );
	
    if (PRINT_RESULTS) $write("Numerator real part: ( ReA * ReB + ImA * ImB ) = %d (%1.8f)\n", NumeR, NumeR/65536.0 );
    if (PRINT_RESULTS) $write("Numerator imag part: ( ReB * ImA - ReA * ImB ) = %d (%1.8f)\n", NumeI, NumeI/65536.0 );
    if (PRINT_RESULTS) $write("Denominator        : ( ReB * ReB + ImB * ImB ) = %d (%1.8f)\n", Denom, Denom/65536.0 );
	
	if ( Denom[31:16] == 16'd0 )
    begin
      if (PRINT_RESULTS) $write("Fixed-point divide error: integer part of denominator is zero\n");
      if (PRINT_RESULTS) $write("This is an overflow condition: the complex quotient does not fit in 16 integer bits\n");
	  // Set final result to unknown:
	  ReY = 32'dx;
      ImY = 32'dx;
    end
	
    if (PRINT_RESULTS) $write("ReY = %d (%1.8f)\n", ReY, ReY/65536.0 );
    if (PRINT_RESULTS) $write("ImY = %d (%1.8f)\n", ImY, ImY/65536.0 );
 	
  end

end
endtask		



//--------------------------------------------------------------------
// Auxiliary functions
//--------------------------------------------------------------------
// Fixed-point multiplication, signed multiplicand and multiplier:
function [31:0] fxpmult (
                          input[15:0] A, 
                          input[15:0] B
						);
reg [15:0] absA;
reg [15:0] absB;
reg [31:0] P;
reg sP;
begin
  sP = A[15] ^ B[15];
  absA = A[15] ? -A : A;
  absB = B[15] ? -B : B;
  P = absA * absB;
  fxpmult = sP ? -P : P;
end
endfunction


//--------------------------------------------------------------------
// Fixed-point division, signed dividend, unsigned divisor:
function [31:0] fxpdiv (
                          input[31:0] A, 
                          input[15:0] B
						);
reg [31:0] absA;
reg sA;
reg [31:0] Q;
begin
  sA = A[31];
  absA = A[31] ? -A : A;
  Q = absA / B;
  fxpdiv = sA ? -Q : Q;
end
endfunction		   

endmodule
